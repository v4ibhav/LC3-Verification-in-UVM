import uvm_pkg::*;
import lc3_test_pkg::*;
module hvl_top();

initial
begin
$display("Entered into hvl top");
run_test();
end

endmodule
