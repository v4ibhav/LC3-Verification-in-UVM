//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
// DESCRIPTION: Protocol specific agent class definition
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
class decode_in_agent  extends uvmf_parameterized_agent #(
                    .CONFIG_T(decode_in_configuration ),
                    .DRIVER_T(decode_in_driver ),
                    .MONITOR_T(decode_in_monitor ),
                    .COVERAGE_T(decode_in_transaction_coverage ),
                    .TRANS_T(decode_in_transaction )
                    );

  `uvm_component_utils( decode_in_agent )

// pragma uvmf custom class_item_additional begin
// pragma uvmf custom class_item_additional end

// ****************************************************************************
// FUNCTION : new()
// This function is the standard SystemVerilog constructor.
//
  function new( string name = "", uvm_component parent = null );
    super.new( name, parent );
  endfunction

// ****************************************************************************
  // FUNCTION: build_phase
  virtual function void build_phase(uvm_phase phase);
// pragma uvmf custom build_phase_pre_super begin
// pragma uvmf custom build_phase_pre_super end
    super.build_phase(phase);
    if (configuration.active_passive == ACTIVE) begin
      // Place sequencer handle into configuration object
      // so that it may be retrieved from configuration 
      // rather than using uvm_config_db
      configuration.sequencer = this.sequencer;
      // configuration.has_coverage = 1;
    end
  endfunction
  
endclass

// pragma uvmf custom external begin
// pragma uvmf custom external end

